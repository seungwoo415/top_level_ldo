VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO strong_arm
  CLASS CORE ;
  ORIGIN 0.43 35.79 ;
  FOREIGN strong_arm -0.43 -35.79 ;
  SIZE 10.32 BY 36.87 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN clock
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 5.875 -5.6 7.455 -5.2 ;
        RECT 2.005 -5.6 3.585 -5.2 ;
      LAYER li1 ;
        RECT 7.225 -2.785 8.255 -2.615 ;
        RECT 8.085 -33.565 8.255 -2.615 ;
        RECT 7.225 -6.025 8.255 -5.855 ;
        RECT 7.225 -33.565 8.255 -33.395 ;
        RECT 7.225 -2.855 7.395 -2.005 ;
        RECT 7.225 -6.025 7.395 -4.705 ;
        RECT 7.225 -34.175 7.395 -33.325 ;
        RECT 2.065 -2.245 7.395 -2.075 ;
        RECT 5.505 -34.105 7.395 -33.935 ;
        RECT 5.505 -2.855 5.675 -2.005 ;
        RECT 5.505 -34.175 5.675 -33.325 ;
        RECT 3.785 -2.855 3.955 -2.005 ;
        RECT 3.785 -34.175 3.955 -33.325 ;
        RECT 2.065 -34.105 3.955 -33.935 ;
        RECT 2.065 -2.855 2.235 -2.005 ;
        RECT 2.065 -6.025 2.235 -4.705 ;
        RECT 2.065 -34.175 2.235 -33.325 ;
        RECT 1.205 -2.785 2.235 -2.615 ;
        RECT 1.205 -6.025 2.235 -5.855 ;
        RECT 1.205 -33.565 2.235 -33.395 ;
        RECT 1.205 -33.565 1.375 -2.615 ;
        RECT 5.505 -5.485 6.105 -5.315 ;
        RECT 5.505 -5.555 5.675 -4.705 ;
        RECT 3.785 -5.555 3.955 -4.705 ;
        RECT 3.355 -5.485 3.955 -5.315 ;
      LAYER mcon ;
        RECT 2.065 -5.485 2.235 -5.315 ;
        RECT 3.355 -5.485 3.525 -5.315 ;
        RECT 5.935 -5.485 6.105 -5.315 ;
        RECT 7.225 -5.485 7.395 -5.315 ;
    END
  END clock
  PIN input_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.505 -25.535 5.675 -24.685 ;
        RECT 3.785 -25.465 5.675 -25.295 ;
        RECT 3.785 -25.535 3.955 -24.685 ;
    END
  END input_n
  PIN input_p
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.865 -25.04 7.025 -24.64 ;
      LAYER li1 ;
        RECT 7.225 -25.535 7.395 -24.685 ;
        RECT 6.795 -24.925 7.395 -24.755 ;
        RECT 2.065 -24.925 3.095 -24.755 ;
        RECT 2.065 -25.535 2.235 -24.685 ;
      LAYER mcon ;
        RECT 2.925 -24.925 3.095 -24.755 ;
        RECT 6.795 -24.925 6.965 -24.755 ;
    END
  END input_p
  PIN output_n
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.18 -9.92 7.44 -0.88 ;
        RECT 5.89 -21.8 6.15 -20.32 ;
        RECT 3.31 -21.8 3.57 -20.32 ;
        RECT 2.02 -9.92 2.28 -0.88 ;
      LAYER met1 ;
        RECT 5.89 -20.72 7.455 -20.32 ;
        RECT 6.305 -9.92 7.455 -9.52 ;
        RECT 7.165 -7.22 7.455 -6.82 ;
        RECT 7.165 -1.28 7.455 -0.88 ;
        RECT 5.445 -21.8 6.15 -21.4 ;
        RECT 3.31 -21.8 4.015 -21.4 ;
        RECT 2.005 -20.72 3.57 -20.32 ;
        RECT 2.005 -9.92 3.155 -9.52 ;
        RECT 2.005 -7.22 2.295 -6.82 ;
        RECT 2.005 -1.28 2.295 -0.88 ;
      LAYER li1 ;
        RECT 7.225 -21.215 7.395 -9.565 ;
        RECT 7.225 -7.715 7.395 -6.325 ;
        RECT 7.225 -1.775 7.395 -0.925 ;
        RECT 5.935 -9.265 6.535 -9.095 ;
        RECT 6.365 -9.805 6.535 -9.095 ;
        RECT 5.505 -8.725 6.105 -8.555 ;
        RECT 5.935 -9.265 6.105 -8.555 ;
        RECT 5.505 -8.795 5.675 -7.945 ;
        RECT 5.505 -22.295 5.675 -21.445 ;
        RECT 3.785 -22.225 5.675 -22.055 ;
        RECT 3.785 -22.295 3.955 -21.445 ;
        RECT 3.785 -8.795 3.955 -7.945 ;
        RECT 3.355 -8.725 3.955 -8.555 ;
        RECT 3.355 -9.265 3.525 -8.555 ;
        RECT 2.925 -9.265 3.525 -9.095 ;
        RECT 2.925 -9.805 3.095 -9.095 ;
        RECT 2.065 -21.215 2.235 -9.565 ;
        RECT 2.065 -7.715 2.235 -6.325 ;
        RECT 2.065 -1.775 2.235 -0.925 ;
      LAYER mcon ;
        RECT 2.065 -1.165 2.235 -0.995 ;
        RECT 2.065 -7.105 2.235 -6.935 ;
        RECT 2.065 -9.805 2.235 -9.635 ;
        RECT 2.065 -20.605 2.235 -20.435 ;
        RECT 2.925 -9.805 3.095 -9.635 ;
        RECT 3.785 -21.685 3.955 -21.515 ;
        RECT 5.505 -21.685 5.675 -21.515 ;
        RECT 6.365 -9.805 6.535 -9.635 ;
        RECT 7.225 -1.165 7.395 -0.995 ;
        RECT 7.225 -7.105 7.395 -6.935 ;
        RECT 7.225 -9.805 7.395 -9.635 ;
        RECT 7.225 -20.605 7.395 -20.435 ;
      LAYER via ;
        RECT 2.075 -1.155 2.225 -1.005 ;
        RECT 2.075 -7.095 2.225 -6.945 ;
        RECT 2.075 -9.795 2.225 -9.645 ;
        RECT 3.365 -20.595 3.515 -20.445 ;
        RECT 3.365 -21.675 3.515 -21.525 ;
        RECT 5.945 -20.595 6.095 -20.445 ;
        RECT 5.945 -21.675 6.095 -21.525 ;
        RECT 7.235 -1.155 7.385 -1.005 ;
        RECT 7.235 -7.095 7.385 -6.945 ;
        RECT 7.235 -9.795 7.385 -9.645 ;
    END
  END output_n
  PIN output_p
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.18 -21.8 7.44 -20.86 ;
        RECT 5.46 -9.38 5.72 -0.88 ;
        RECT 3.74 -9.38 4 -0.88 ;
        RECT 2.02 -21.8 2.28 -20.86 ;
      LAYER met1 ;
        RECT 7.165 -21.8 7.455 -21.4 ;
        RECT 5.445 -9.38 7.455 -8.98 ;
        RECT 2.02 -21.26 7.44 -20.86 ;
        RECT 5.445 -6.68 5.735 -6.28 ;
        RECT 5.445 -1.28 5.735 -0.88 ;
        RECT 2.005 -9.38 4.015 -8.98 ;
        RECT 3.725 -6.68 4.015 -6.28 ;
        RECT 3.725 -1.28 4.015 -0.88 ;
        RECT 2.005 -21.8 2.295 -21.4 ;
      LAYER li1 ;
        RECT 7.225 -22.295 7.395 -21.445 ;
        RECT 7.225 -9.265 7.395 -7.945 ;
        RECT 5.505 -21.215 5.675 -9.095 ;
        RECT 5.505 -7.715 5.675 -6.325 ;
        RECT 5.505 -1.775 5.675 -0.925 ;
        RECT 3.785 -21.215 3.955 -9.095 ;
        RECT 3.785 -7.715 3.955 -6.325 ;
        RECT 3.785 -1.775 3.955 -0.925 ;
        RECT 2.065 -22.295 2.235 -21.445 ;
        RECT 2.065 -9.265 2.235 -7.945 ;
      LAYER mcon ;
        RECT 2.065 -9.265 2.235 -9.095 ;
        RECT 2.065 -21.685 2.235 -21.515 ;
        RECT 3.785 -1.165 3.955 -0.995 ;
        RECT 3.785 -6.565 3.955 -6.395 ;
        RECT 3.785 -9.265 3.955 -9.095 ;
        RECT 3.785 -21.145 3.955 -20.975 ;
        RECT 5.505 -1.165 5.675 -0.995 ;
        RECT 5.505 -6.565 5.675 -6.395 ;
        RECT 5.505 -9.265 5.675 -9.095 ;
        RECT 5.505 -21.145 5.675 -20.975 ;
        RECT 7.225 -9.265 7.395 -9.095 ;
        RECT 7.225 -21.685 7.395 -21.515 ;
      LAYER via ;
        RECT 2.075 -21.135 2.225 -20.985 ;
        RECT 2.075 -21.675 2.225 -21.525 ;
        RECT 3.795 -1.155 3.945 -1.005 ;
        RECT 3.795 -6.555 3.945 -6.405 ;
        RECT 3.795 -9.255 3.945 -9.105 ;
        RECT 5.515 -1.155 5.665 -1.005 ;
        RECT 5.515 -6.555 5.665 -6.405 ;
        RECT 5.515 -9.255 5.665 -9.105 ;
        RECT 7.235 -21.135 7.385 -20.985 ;
        RECT 7.235 -21.675 7.385 -21.525 ;
    END
  END output_p
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 5.015 -7.76 9.605 -7.36 ;
        RECT 5.015 -4.52 9.605 -4.12 ;
        RECT 8.455 -1.82 9.605 -1.42 ;
        RECT 6.735 -1.82 7.885 -1.42 ;
        RECT 5.015 -1.82 6.165 -1.42 ;
        RECT -0.145 -7.76 4.445 -7.36 ;
        RECT -0.145 -4.52 4.445 -4.12 ;
        RECT 3.295 -1.82 4.445 -1.42 ;
        RECT 1.575 -1.82 2.725 -1.42 ;
        RECT -0.145 -1.82 1.005 -1.42 ;
      LAYER li1 ;
        RECT 4.995 -0.085 9.625 0.625 ;
        RECT 9.375 -1.775 9.545 0.625 ;
        RECT 6.795 -1.775 6.965 0.625 ;
        RECT 5.075 -1.775 5.245 0.625 ;
        RECT 9.375 -7.715 9.545 -6.325 ;
        RECT 9.375 -4.475 9.545 -3.625 ;
        RECT 8.945 -3.865 9.545 -3.695 ;
        RECT 8.945 -8.795 9.115 -0.925 ;
        RECT 8.515 -7.715 8.685 -6.325 ;
        RECT 8.515 -4.475 8.685 -3.625 ;
        RECT 8.515 -1.775 8.685 -0.925 ;
        RECT 7.655 -7.715 7.825 -6.325 ;
        RECT 7.655 -4.475 7.825 -3.625 ;
        RECT 7.655 -1.775 7.825 -0.925 ;
        RECT 6.795 -7.715 6.965 -6.325 ;
        RECT 6.795 -4.475 6.965 -3.625 ;
        RECT 5.935 -7.715 6.105 -6.325 ;
        RECT 5.935 -4.475 6.105 -3.625 ;
        RECT 5.935 -1.775 6.105 -0.925 ;
        RECT 5.075 -7.715 5.245 -6.325 ;
        RECT 4.215 -7.645 5.245 -7.475 ;
        RECT 4.215 -7.715 4.385 -6.325 ;
        RECT 5.075 -4.475 5.245 -3.625 ;
        RECT -0.165 -0.085 4.465 0.625 ;
        RECT 4.215 -1.775 4.385 0.625 ;
        RECT 2.495 -1.775 2.665 0.625 ;
        RECT -0.085 -1.775 0.085 0.625 ;
        RECT 4.215 -4.475 4.385 -3.625 ;
        RECT 3.355 -7.715 3.525 -6.325 ;
        RECT 3.355 -4.475 3.525 -3.625 ;
        RECT 3.355 -1.775 3.525 -0.925 ;
        RECT 2.495 -7.715 2.665 -6.325 ;
        RECT 2.495 -4.475 2.665 -3.625 ;
        RECT 1.635 -7.715 1.805 -6.325 ;
        RECT 1.635 -4.475 1.805 -3.625 ;
        RECT 1.635 -1.775 1.805 -0.925 ;
        RECT 0.775 -7.715 0.945 -6.325 ;
        RECT 0.775 -4.475 0.945 -3.625 ;
        RECT 0.775 -1.775 0.945 -0.925 ;
        RECT 0.345 -8.795 0.515 -0.925 ;
        RECT -0.085 -3.865 0.515 -3.695 ;
        RECT -0.085 -4.475 0.085 -3.625 ;
        RECT -0.085 -7.715 0.085 -6.325 ;
      LAYER mcon ;
        RECT -0.085 -1.705 0.085 -1.535 ;
        RECT -0.085 -4.405 0.085 -4.235 ;
        RECT -0.085 -7.645 0.085 -7.475 ;
        RECT 0.345 -1.705 0.515 -1.535 ;
        RECT 0.345 -7.645 0.515 -7.475 ;
        RECT 0.775 -1.705 0.945 -1.535 ;
        RECT 0.775 -4.405 0.945 -4.235 ;
        RECT 0.775 -7.645 0.945 -7.475 ;
        RECT 1.635 -1.705 1.805 -1.535 ;
        RECT 1.635 -4.405 1.805 -4.235 ;
        RECT 1.635 -7.645 1.805 -7.475 ;
        RECT 2.495 -1.705 2.665 -1.535 ;
        RECT 2.495 -4.405 2.665 -4.235 ;
        RECT 2.495 -7.645 2.665 -7.475 ;
        RECT 3.355 -1.705 3.525 -1.535 ;
        RECT 3.355 -4.405 3.525 -4.235 ;
        RECT 3.355 -7.645 3.525 -7.475 ;
        RECT 4.215 -1.705 4.385 -1.535 ;
        RECT 4.215 -4.405 4.385 -4.235 ;
        RECT 4.215 -7.645 4.385 -7.475 ;
        RECT 5.075 -1.705 5.245 -1.535 ;
        RECT 5.075 -4.405 5.245 -4.235 ;
        RECT 5.075 -7.645 5.245 -7.475 ;
        RECT 5.935 -1.705 6.105 -1.535 ;
        RECT 5.935 -4.405 6.105 -4.235 ;
        RECT 5.935 -7.645 6.105 -7.475 ;
        RECT 6.795 -1.705 6.965 -1.535 ;
        RECT 6.795 -4.405 6.965 -4.235 ;
        RECT 6.795 -7.645 6.965 -7.475 ;
        RECT 7.655 -1.705 7.825 -1.535 ;
        RECT 7.655 -4.405 7.825 -4.235 ;
        RECT 7.655 -7.645 7.825 -7.475 ;
        RECT 8.515 -1.705 8.685 -1.535 ;
        RECT 8.515 -4.405 8.685 -4.235 ;
        RECT 8.515 -7.645 8.685 -7.475 ;
        RECT 8.945 -1.705 9.115 -1.535 ;
        RECT 8.945 -7.645 9.115 -7.475 ;
        RECT 9.375 -1.705 9.545 -1.535 ;
        RECT 9.375 -4.405 9.545 -4.235 ;
        RECT 9.375 -7.645 9.545 -7.475 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 6.735 -28.28 9.605 -27.88 ;
        RECT 8.455 -24.5 9.605 -24.1 ;
        RECT 8.455 -18.02 9.605 -17.62 ;
        RECT 3.295 -28.28 6.165 -27.88 ;
        RECT -0.145 -28.28 2.725 -27.88 ;
        RECT -0.145 -24.5 1.005 -24.1 ;
        RECT -0.145 -18.02 1.005 -17.62 ;
      LAYER li1 ;
        RECT 4.995 -35.725 9.625 -35.015 ;
        RECT 9.375 -33.095 9.545 -26.305 ;
        RECT 8.945 -26.545 9.545 -26.375 ;
        RECT 8.945 -35.725 9.115 -9.565 ;
        RECT 8.515 -18.985 9.115 -18.815 ;
        RECT 8.515 -21.215 8.685 -9.565 ;
        RECT 9.375 -24.455 9.545 -23.065 ;
        RECT 9.375 -21.215 9.545 -9.565 ;
        RECT 8.515 -33.095 8.685 -26.305 ;
        RECT 8.515 -24.455 8.685 -23.065 ;
        RECT 7.655 -33.095 7.825 -26.305 ;
        RECT 6.795 -33.095 6.965 -26.305 ;
        RECT 5.935 -27.625 6.965 -27.455 ;
        RECT 5.935 -33.095 6.105 -26.305 ;
        RECT 5.075 -33.095 5.245 -26.305 ;
        RECT -0.165 -35.725 4.465 -35.015 ;
        RECT 0.775 -21.215 0.945 -9.565 ;
        RECT 0.345 -18.985 0.945 -18.815 ;
        RECT 0.345 -35.725 0.515 -9.565 ;
        RECT -0.085 -26.545 0.515 -26.375 ;
        RECT -0.085 -33.095 0.085 -26.305 ;
        RECT 4.215 -33.095 4.385 -26.305 ;
        RECT 3.355 -33.095 3.525 -26.305 ;
        RECT 2.495 -27.625 3.525 -27.455 ;
        RECT 2.495 -33.095 2.665 -26.305 ;
        RECT 1.635 -33.095 1.805 -26.305 ;
        RECT 0.775 -33.095 0.945 -26.305 ;
        RECT 0.775 -24.455 0.945 -23.065 ;
        RECT -0.085 -24.455 0.085 -23.065 ;
        RECT -0.085 -21.215 0.085 -9.565 ;
      LAYER mcon ;
        RECT -0.085 -17.905 0.085 -17.735 ;
        RECT -0.085 -24.385 0.085 -24.215 ;
        RECT -0.085 -28.165 0.085 -27.995 ;
        RECT 0.345 -24.385 0.515 -24.215 ;
        RECT 0.775 -17.905 0.945 -17.735 ;
        RECT 0.775 -24.385 0.945 -24.215 ;
        RECT 0.775 -28.165 0.945 -27.995 ;
        RECT 1.635 -28.165 1.805 -27.995 ;
        RECT 2.495 -28.165 2.665 -27.995 ;
        RECT 3.355 -28.165 3.525 -27.995 ;
        RECT 4.215 -28.165 4.385 -27.995 ;
        RECT 5.075 -28.165 5.245 -27.995 ;
        RECT 5.935 -28.165 6.105 -27.995 ;
        RECT 6.795 -28.165 6.965 -27.995 ;
        RECT 7.655 -28.165 7.825 -27.995 ;
        RECT 8.515 -17.905 8.685 -17.735 ;
        RECT 8.515 -24.385 8.685 -24.215 ;
        RECT 8.515 -28.165 8.685 -27.995 ;
        RECT 8.945 -24.385 9.115 -24.215 ;
        RECT 9.375 -17.905 9.545 -17.735 ;
        RECT 9.375 -24.385 9.545 -24.215 ;
        RECT 9.375 -28.165 9.545 -27.995 ;
    END
  END vss
  OBS
    LAYER mcon ;
      RECT 7.655 -24.385 7.825 -24.215 ;
      RECT 7.655 -17.905 7.825 -17.735 ;
      RECT 6.795 -24.385 6.965 -24.215 ;
      RECT 6.795 -17.905 6.965 -17.735 ;
      RECT 5.935 -24.385 6.105 -24.215 ;
      RECT 5.935 -17.905 6.105 -17.735 ;
      RECT 5.505 -3.865 5.675 -3.695 ;
      RECT 5.075 -24.385 5.245 -24.215 ;
      RECT 5.075 -17.905 5.245 -17.735 ;
      RECT 5.075 -9.265 5.245 -9.095 ;
      RECT 4.215 -24.385 4.385 -24.215 ;
      RECT 4.215 -17.905 4.385 -17.735 ;
      RECT 4.215 -9.265 4.385 -9.095 ;
      RECT 3.785 -3.865 3.955 -3.695 ;
      RECT 3.355 -24.385 3.525 -24.215 ;
      RECT 3.355 -17.905 3.525 -17.735 ;
      RECT 2.495 -24.385 2.665 -24.215 ;
      RECT 2.495 -17.905 2.665 -17.735 ;
      RECT 1.635 -24.385 1.805 -24.215 ;
      RECT 1.635 -17.905 1.805 -17.735 ;
    LAYER met1 ;
      RECT 6.735 -24.5 7.885 -24.1 ;
      RECT 6.735 -18.02 7.885 -17.62 ;
      RECT 5.015 -24.5 6.165 -24.1 ;
      RECT 5.015 -18.02 6.165 -17.62 ;
      RECT 5.03 -3.98 5.735 -3.58 ;
      RECT 5.015 -9.38 5.305 -8.98 ;
      RECT 3.295 -24.5 4.445 -24.1 ;
      RECT 3.295 -18.02 4.445 -17.62 ;
      RECT 4.155 -9.38 4.445 -8.98 ;
      RECT 3.725 -3.98 4.43 -3.58 ;
      RECT 1.575 -24.5 2.725 -24.1 ;
      RECT 1.575 -18.02 2.725 -17.62 ;
    LAYER via ;
      RECT 5.085 -9.255 5.235 -9.105 ;
      RECT 5.085 -3.855 5.235 -3.705 ;
      RECT 4.225 -9.255 4.375 -9.105 ;
      RECT 4.225 -3.855 4.375 -3.705 ;
    LAYER met2 ;
      RECT 5.03 -9.38 5.29 -3.58 ;
      RECT 4.17 -9.38 4.43 -3.58 ;
    LAYER li1 ;
      RECT 6.795 -24.455 6.965 -23.065 ;
      RECT 5.935 -26.005 6.105 -23.065 ;
      RECT 5.935 -23.845 6.965 -23.675 ;
      RECT 5.505 -26.005 7.395 -25.835 ;
      RECT 7.225 -33.095 7.395 -25.835 ;
      RECT 5.505 -33.095 5.675 -25.835 ;
      RECT 6.365 -3.325 7.395 -3.155 ;
      RECT 7.225 -4.475 7.395 -3.155 ;
      RECT 2.065 -3.325 3.095 -3.155 ;
      RECT 2.925 -8.725 3.095 -3.155 ;
      RECT 6.365 -8.725 6.535 -3.155 ;
      RECT 2.065 -4.475 2.235 -3.155 ;
      RECT 2.925 -6.025 6.535 -5.855 ;
      RECT 6.365 -8.725 6.965 -8.555 ;
      RECT 6.795 -22.765 6.965 -8.555 ;
      RECT 2.495 -8.725 3.095 -8.555 ;
      RECT 2.495 -22.765 2.665 -8.555 ;
      RECT 6.795 -22.765 7.395 -22.595 ;
      RECT 7.225 -24.455 7.395 -22.595 ;
      RECT 2.065 -22.765 2.665 -22.595 ;
      RECT 2.065 -24.455 2.235 -22.595 ;
      RECT 5.935 -22.765 6.105 -9.565 ;
      RECT 5.505 -22.765 6.105 -22.595 ;
      RECT 5.505 -24.455 5.675 -22.595 ;
      RECT 5.075 -24.455 5.245 -23.065 ;
      RECT 4.215 -24.455 4.385 -23.065 ;
      RECT 4.215 -24.385 5.245 -24.215 ;
      RECT 3.355 -26.005 3.525 -23.065 ;
      RECT 2.495 -24.455 2.665 -23.065 ;
      RECT 2.495 -23.845 3.525 -23.675 ;
      RECT 2.065 -26.005 3.955 -25.835 ;
      RECT 3.785 -33.095 3.955 -25.835 ;
      RECT 2.065 -33.095 2.235 -25.835 ;
      RECT 3.355 -22.765 3.525 -9.565 ;
      RECT 3.355 -22.765 3.955 -22.595 ;
      RECT 3.785 -24.455 3.955 -22.595 ;
      RECT 7.655 -24.455 7.825 -23.065 ;
      RECT 7.655 -21.215 7.825 -9.565 ;
      RECT 5.505 -4.475 5.675 -3.625 ;
      RECT 5.075 -21.215 5.245 -9.095 ;
      RECT 4.215 -21.215 4.385 -9.095 ;
      RECT 3.785 -4.475 3.955 -3.625 ;
      RECT 1.635 -24.455 1.805 -23.065 ;
      RECT 1.635 -21.215 1.805 -9.565 ;
  END
END strong_arm

END LIBRARY
