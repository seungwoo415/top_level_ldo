VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO pass_transistors
  CLASS CORE ;
  ORIGIN -0.305 9.87 ;
  FOREIGN pass_transistors 0.305 -9.87 ;
  SIZE 22.775 BY 24.16 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.305 -0.56 0.665 12.865 ;
        RECT 0.355 -0.56 0.615 12.93 ;
      LAYER li1 ;
        RECT 20.935 -0.17 21.465 0.16 ;
        RECT 20.89 12.38 21.42 12.71 ;
        RECT 19.88 -1.87 20.05 -0.095 ;
        RECT 19.865 10.48 20.035 12.245 ;
        RECT 18.825 -1.87 18.995 -0.095 ;
        RECT 18.805 10.48 18.975 12.26 ;
        RECT 17.765 -1.87 17.935 -0.095 ;
        RECT 17.745 10.48 17.915 12.24 ;
        RECT 17.215 -1.6 17.385 -0.91 ;
        RECT 17.085 10.78 17.255 11.47 ;
        RECT 16.09 -1.87 16.26 -0.095 ;
        RECT 15.88 10.48 16.05 12.24 ;
        RECT 15.03 -1.87 15.2 -0.095 ;
        RECT 14.82 10.48 14.99 12.23 ;
        RECT 13.97 -1.865 14.14 -0.09 ;
        RECT 13.77 10.485 13.94 12.24 ;
        RECT 12.91 -1.865 13.08 -0.09 ;
        RECT 12.715 10.485 12.885 12.24 ;
        RECT 11.855 -1.865 12.025 -0.09 ;
        RECT 11.66 10.485 11.83 12.24 ;
        RECT 10.8 -1.865 10.97 -0.09 ;
        RECT 10.6 10.485 10.77 12.24 ;
        RECT 10.305 -1.595 10.475 -0.905 ;
        RECT 9.935 10.72 10.105 11.41 ;
        RECT 9.185 -1.865 9.355 -0.085 ;
        RECT 8.745 10.485 8.915 12.25 ;
        RECT 8.125 -1.865 8.295 -0.09 ;
        RECT 7.69 10.485 7.86 12.25 ;
        RECT 7.065 -1.865 7.235 -0.09 ;
        RECT 6.635 10.485 6.805 12.245 ;
        RECT 6.005 -1.865 6.175 -0.09 ;
        RECT 5.575 10.485 5.745 12.245 ;
        RECT 4.95 -1.865 5.12 -0.09 ;
        RECT 4.515 10.485 4.685 12.23 ;
        RECT 3.89 -1.865 4.06 -0.09 ;
        RECT 3.455 10.485 3.625 12.23 ;
        RECT 2.83 -1.865 3 -0.09 ;
        RECT 2.395 10.485 2.565 12.225 ;
        RECT 1.91 0.03 2.44 0.36 ;
        RECT 1.515 12.395 2.045 12.725 ;
      LAYER met1 ;
        RECT 0.335 12.395 22.415 12.935 ;
        RECT 19.835 11.935 20.065 12.935 ;
        RECT 18.775 11.95 19.005 12.935 ;
        RECT 17.715 11.93 17.945 12.935 ;
        RECT 17.055 10.8 17.285 12.935 ;
        RECT 15.85 11.93 16.08 12.935 ;
        RECT 14.79 11.92 15.02 12.935 ;
        RECT 13.74 11.93 13.97 12.935 ;
        RECT 12.685 11.93 12.915 12.935 ;
        RECT 11.63 11.93 11.86 12.935 ;
        RECT 10.57 11.93 10.8 12.935 ;
        RECT 9.905 10.74 10.135 12.935 ;
        RECT 8.715 11.94 8.945 12.935 ;
        RECT 7.66 11.94 7.89 12.935 ;
        RECT 6.605 11.935 6.835 12.935 ;
        RECT 5.545 11.935 5.775 12.935 ;
        RECT 4.485 11.92 4.715 12.935 ;
        RECT 3.425 11.92 3.655 12.935 ;
        RECT 2.365 11.915 2.595 12.935 ;
        RECT 0.355 12.29 0.615 12.935 ;
        RECT 0.315 0.045 22.33 0.585 ;
        RECT 20.905 -0.15 21.495 0.585 ;
        RECT 19.85 -0.405 20.08 0.585 ;
        RECT 18.795 -0.405 19.025 0.585 ;
        RECT 17.735 -0.405 17.965 0.585 ;
        RECT 17.185 -1.58 17.415 0.585 ;
        RECT 16.06 -0.405 16.29 0.585 ;
        RECT 15 -0.405 15.23 0.585 ;
        RECT 13.94 -0.4 14.17 0.585 ;
        RECT 12.88 -0.4 13.11 0.585 ;
        RECT 11.825 -0.4 12.055 0.585 ;
        RECT 10.77 -0.4 11 0.585 ;
        RECT 10.275 -1.575 10.505 0.585 ;
        RECT 9.155 -0.395 9.385 0.585 ;
        RECT 8.095 -0.4 8.325 0.585 ;
        RECT 7.035 -0.4 7.265 0.585 ;
        RECT 5.975 -0.4 6.205 0.585 ;
        RECT 4.92 -0.4 5.15 0.585 ;
        RECT 3.86 -0.4 4.09 0.585 ;
        RECT 2.8 -0.4 3.03 0.585 ;
        RECT 0.36 -0.035 0.62 0.605 ;
      LAYER mcon ;
        RECT 1.515 12.475 1.685 12.645 ;
        RECT 1.875 12.475 2.045 12.645 ;
        RECT 1.91 0.11 2.08 0.28 ;
        RECT 2.27 0.11 2.44 0.28 ;
        RECT 2.395 11.975 2.565 12.145 ;
        RECT 2.83 -0.34 3 -0.17 ;
        RECT 3.455 11.98 3.625 12.15 ;
        RECT 3.89 -0.34 4.06 -0.17 ;
        RECT 4.515 11.98 4.685 12.15 ;
        RECT 4.95 -0.34 5.12 -0.17 ;
        RECT 5.575 11.995 5.745 12.165 ;
        RECT 6.005 -0.34 6.175 -0.17 ;
        RECT 6.635 11.995 6.805 12.165 ;
        RECT 7.065 -0.34 7.235 -0.17 ;
        RECT 7.69 12 7.86 12.17 ;
        RECT 8.125 -0.34 8.295 -0.17 ;
        RECT 8.745 12 8.915 12.17 ;
        RECT 9.185 -0.335 9.355 -0.165 ;
        RECT 9.935 11.16 10.105 11.33 ;
        RECT 9.935 10.8 10.105 10.97 ;
        RECT 10.305 -1.155 10.475 -0.985 ;
        RECT 10.305 -1.515 10.475 -1.345 ;
        RECT 10.6 11.99 10.77 12.16 ;
        RECT 10.8 -0.34 10.97 -0.17 ;
        RECT 11.66 11.99 11.83 12.16 ;
        RECT 11.855 -0.34 12.025 -0.17 ;
        RECT 12.715 11.99 12.885 12.16 ;
        RECT 12.91 -0.34 13.08 -0.17 ;
        RECT 13.77 11.99 13.94 12.16 ;
        RECT 13.97 -0.34 14.14 -0.17 ;
        RECT 14.82 11.98 14.99 12.15 ;
        RECT 15.03 -0.345 15.2 -0.175 ;
        RECT 15.88 11.99 16.05 12.16 ;
        RECT 16.09 -0.345 16.26 -0.175 ;
        RECT 17.085 11.22 17.255 11.39 ;
        RECT 17.085 10.86 17.255 11.03 ;
        RECT 17.215 -1.16 17.385 -0.99 ;
        RECT 17.215 -1.52 17.385 -1.35 ;
        RECT 17.745 11.99 17.915 12.16 ;
        RECT 17.765 -0.345 17.935 -0.175 ;
        RECT 18.805 12.01 18.975 12.18 ;
        RECT 18.825 -0.345 18.995 -0.175 ;
        RECT 19.865 11.995 20.035 12.165 ;
        RECT 19.88 -0.345 20.05 -0.175 ;
        RECT 20.89 12.46 21.06 12.63 ;
        RECT 20.935 -0.09 21.105 0.08 ;
        RECT 21.25 12.46 21.42 12.63 ;
        RECT 21.295 -0.09 21.465 0.08 ;
      LAYER via ;
        RECT 0.41 12.695 0.56 12.845 ;
        RECT 0.41 12.375 0.56 12.525 ;
        RECT 0.415 0.37 0.565 0.52 ;
        RECT 0.415 0.05 0.565 0.2 ;
    END
  END VDD
  PIN Vg_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095 -2.46 3.265 -2.13 ;
      LAYER met1 ;
        RECT 2.805 -2.44 3.295 -2.15 ;
      LAYER mcon ;
        RECT 3.095 -2.38 3.265 -2.21 ;
    END
  END Vg_0
  PIN Vg_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.155 -2.895 4.325 -2.11 ;
      LAYER met1 ;
        RECT 2.81 -2.875 4.355 -2.585 ;
        RECT 4.02 -2.42 4.355 -2.13 ;
      LAYER mcon ;
        RECT 4.155 -2.36 4.325 -2.19 ;
        RECT 4.155 -2.815 4.325 -2.645 ;
    END
  END Vg_1
  PIN Vg_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.235 -7.22 14.405 -2.1 ;
      LAYER met1 ;
        RECT 3.5 -7.2 14.435 -6.91 ;
        RECT 13.975 -2.41 14.435 -2.12 ;
      LAYER mcon ;
        RECT 14.235 -2.35 14.405 -2.18 ;
        RECT 14.235 -7.14 14.405 -6.97 ;
    END
  END Vg_10
  PIN Vg_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.295 -7.76 15.465 -2.11 ;
      LAYER met1 ;
        RECT 3.535 -7.74 15.495 -7.45 ;
        RECT 15.005 -2.42 15.495 -2.13 ;
      LAYER mcon ;
        RECT 15.295 -2.36 15.465 -2.19 ;
        RECT 15.295 -7.68 15.465 -7.51 ;
    END
  END Vg_11
  PIN Vg_12
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.36 -8.325 16.53 -2.105 ;
      LAYER met1 ;
        RECT 3.59 -8.305 16.56 -8.015 ;
        RECT 16.15 -2.415 16.56 -2.125 ;
      LAYER mcon ;
        RECT 16.36 -2.355 16.53 -2.185 ;
        RECT 16.36 -8.245 16.53 -8.075 ;
    END
  END Vg_12
  PIN Vg_13
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.03 -8.905 18.2 -2.13 ;
      LAYER met1 ;
        RECT 3.735 -8.885 18.23 -8.595 ;
        RECT 17.825 -2.44 18.23 -2.15 ;
      LAYER mcon ;
        RECT 18.03 -2.38 18.2 -2.21 ;
        RECT 18.03 -8.825 18.2 -8.655 ;
    END
  END Vg_13
  PIN Vg_14
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.09 -9.4 19.26 -2.12 ;
      LAYER met1 ;
        RECT 3.8 -9.38 19.29 -9.09 ;
        RECT 18.845 -2.43 19.29 -2.14 ;
      LAYER mcon ;
        RECT 19.09 -2.37 19.26 -2.2 ;
        RECT 19.09 -9.32 19.26 -9.15 ;
    END
  END Vg_14
  PIN Vg_15
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 20.15 -9.87 20.32 -2.125 ;
      LAYER met1 ;
        RECT 3.85 -9.85 20.35 -9.56 ;
        RECT 19.905 -2.435 20.35 -2.145 ;
      LAYER mcon ;
        RECT 20.15 -2.375 20.32 -2.205 ;
        RECT 20.15 -9.79 20.32 -9.62 ;
    END
  END Vg_15
  PIN Vg_16
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.66 9.895 2.83 10.225 ;
      LAYER met1 ;
        RECT 2.34 9.915 2.86 10.205 ;
      LAYER mcon ;
        RECT 2.66 9.975 2.83 10.145 ;
    END
  END Vg_16
  PIN Vg_17
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.715 9.435 3.885 10.215 ;
      LAYER met1 ;
        RECT 2.49 9.455 3.915 9.745 ;
        RECT 3.5 9.905 3.915 10.195 ;
      LAYER mcon ;
        RECT 3.715 9.965 3.885 10.135 ;
        RECT 3.715 9.515 3.885 9.685 ;
    END
  END Vg_17
  PIN Vg_18
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.775 8.975 4.945 10.225 ;
      LAYER met1 ;
        RECT 2.545 8.995 4.975 9.285 ;
        RECT 4.51 9.915 4.975 10.205 ;
      LAYER mcon ;
        RECT 4.775 9.975 4.945 10.145 ;
        RECT 4.775 9.055 4.945 9.225 ;
    END
  END Vg_18
  PIN Vg_19
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.845 8.52 6.015 10.23 ;
      LAYER met1 ;
        RECT 2.61 8.54 6.045 8.83 ;
        RECT 5.625 9.92 6.045 10.21 ;
      LAYER mcon ;
        RECT 5.845 9.98 6.015 10.15 ;
        RECT 5.845 8.6 6.015 8.77 ;
    END
  END Vg_19
  PIN Vg_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.22 -3.34 5.39 -2.1 ;
      LAYER met1 ;
        RECT 2.99 -3.32 5.42 -3.03 ;
        RECT 5.02 -2.41 5.42 -2.12 ;
      LAYER mcon ;
        RECT 5.22 -2.35 5.39 -2.18 ;
        RECT 5.22 -3.26 5.39 -3.09 ;
    END
  END Vg_2
  PIN Vg_20
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.9 8.07 7.07 10.235 ;
      LAYER met1 ;
        RECT 2.665 8.09 7.1 8.38 ;
        RECT 6.745 9.925 7.1 10.215 ;
      LAYER mcon ;
        RECT 6.9 9.985 7.07 10.155 ;
        RECT 6.9 8.15 7.07 8.32 ;
    END
  END Vg_20
  PIN Vg_21
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.96 7.595 8.13 10.235 ;
      LAYER met1 ;
        RECT 2.725 7.615 8.16 7.905 ;
        RECT 7.825 9.925 8.16 10.215 ;
      LAYER mcon ;
        RECT 7.96 9.985 8.13 10.155 ;
        RECT 7.96 7.675 8.13 7.845 ;
    END
  END Vg_21
  PIN Vg_22
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.015 7.135 9.185 10.235 ;
      LAYER met1 ;
        RECT 2.785 7.155 9.215 7.445 ;
        RECT 8.85 9.925 9.215 10.215 ;
      LAYER mcon ;
        RECT 9.015 9.985 9.185 10.155 ;
        RECT 9.015 7.215 9.185 7.385 ;
    END
  END Vg_22
  PIN Vg_23
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.865 6.64 11.035 10.23 ;
      LAYER met1 ;
        RECT 3.125 6.66 11.065 6.95 ;
        RECT 10.655 9.92 11.065 10.21 ;
      LAYER mcon ;
        RECT 10.865 9.98 11.035 10.15 ;
        RECT 10.865 6.72 11.035 6.89 ;
    END
  END Vg_23
  PIN Vg_24
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.925 6.12 12.095 10.24 ;
      LAYER met1 ;
        RECT 3.19 6.14 12.125 6.43 ;
        RECT 11.665 9.93 12.125 10.22 ;
      LAYER mcon ;
        RECT 11.925 9.99 12.095 10.16 ;
        RECT 11.925 6.2 12.095 6.37 ;
    END
  END Vg_24
  PIN Vg_25
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.985 5.57 13.155 10.24 ;
      LAYER met1 ;
        RECT 3.25 5.59 13.185 5.88 ;
        RECT 12.77 9.93 13.185 10.22 ;
      LAYER mcon ;
        RECT 12.985 9.99 13.155 10.16 ;
        RECT 12.985 5.65 13.155 5.82 ;
    END
  END Vg_25
  PIN Vg_26
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.04 5.13 14.21 10.255 ;
      LAYER met1 ;
        RECT 3.305 5.15 14.24 5.44 ;
        RECT 13.79 9.945 14.24 10.235 ;
      LAYER mcon ;
        RECT 14.04 10.005 14.21 10.175 ;
        RECT 14.04 5.21 14.21 5.38 ;
    END
  END Vg_26
  PIN Vg_27
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.09 4.59 15.26 10.245 ;
      LAYER met1 ;
        RECT 3.33 4.61 15.29 4.9 ;
        RECT 14.92 9.935 15.29 10.225 ;
      LAYER mcon ;
        RECT 15.09 9.995 15.26 10.165 ;
        RECT 15.09 4.67 15.26 4.84 ;
    END
  END Vg_27
  PIN Vg_28
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.145 4.02 16.315 10.245 ;
      LAYER met1 ;
        RECT 3.375 4.04 16.345 4.33 ;
        RECT 15.965 9.935 16.345 10.225 ;
      LAYER mcon ;
        RECT 16.145 9.995 16.315 10.165 ;
        RECT 16.145 4.1 16.315 4.27 ;
    END
  END Vg_28
  PIN Vg_29
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.015 3.485 18.185 10.255 ;
      LAYER met1 ;
        RECT 3.72 3.505 18.215 3.795 ;
        RECT 17.84 9.945 18.215 10.235 ;
      LAYER mcon ;
        RECT 18.015 10.005 18.185 10.175 ;
        RECT 18.015 3.565 18.185 3.735 ;
    END
  END Vg_29
  PIN Vg_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.27 -3.825 6.44 -2.105 ;
      LAYER met1 ;
        RECT 3.035 -3.805 6.47 -3.515 ;
        RECT 6.065 -2.415 6.47 -2.125 ;
      LAYER mcon ;
        RECT 6.27 -2.355 6.44 -2.185 ;
        RECT 6.27 -3.745 6.44 -3.575 ;
    END
  END Vg_3
  PIN Vg_30
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.07 2.995 19.24 10.245 ;
      LAYER met1 ;
        RECT 3.775 3.015 19.27 3.305 ;
        RECT 18.895 9.935 19.27 10.225 ;
      LAYER mcon ;
        RECT 19.07 9.995 19.24 10.165 ;
        RECT 19.07 3.075 19.24 3.245 ;
    END
  END Vg_30
  PIN Vg_31
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 20.135 2.52 20.305 10.245 ;
      LAYER met1 ;
        RECT 3.835 2.54 20.335 2.83 ;
        RECT 19.91 9.935 20.335 10.225 ;
      LAYER mcon ;
        RECT 20.135 9.995 20.305 10.165 ;
        RECT 20.135 2.6 20.305 2.77 ;
    END
  END Vg_31
  PIN Vg_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.33 -4.27 7.5 -2.11 ;
      LAYER met1 ;
        RECT 3.095 -4.25 7.53 -3.96 ;
        RECT 7.125 -2.415 7.53 -2.13 ;
        RECT 7.3 -2.42 7.53 -2.13 ;
      LAYER mcon ;
        RECT 7.33 -2.36 7.5 -2.19 ;
        RECT 7.33 -4.19 7.5 -4.02 ;
    END
  END Vg_4
  PIN Vg_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.395 -4.74 8.565 -2.11 ;
      LAYER met1 ;
        RECT 3.16 -4.72 8.595 -4.43 ;
        RECT 8.22 -2.42 8.595 -2.13 ;
      LAYER mcon ;
        RECT 8.395 -2.36 8.565 -2.19 ;
        RECT 8.395 -4.66 8.565 -4.49 ;
    END
  END Vg_5
  PIN Vg_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.455 -5.215 9.625 -2.12 ;
      LAYER met1 ;
        RECT 3.225 -5.195 9.655 -4.905 ;
        RECT 9.265 -2.43 9.655 -2.14 ;
        RECT 9.265 -2.43 9.425 -2.135 ;
      LAYER mcon ;
        RECT 9.455 -2.37 9.625 -2.2 ;
        RECT 9.455 -5.135 9.625 -4.965 ;
    END
  END Vg_6
  PIN Vg_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.07 -5.71 11.24 -2.12 ;
      LAYER met1 ;
        RECT 3.33 -5.69 11.27 -5.4 ;
        RECT 10.9 -2.43 11.27 -2.14 ;
      LAYER mcon ;
        RECT 11.07 -2.37 11.24 -2.2 ;
        RECT 11.07 -5.63 11.24 -5.46 ;
    END
  END Vg_7
  PIN Vg_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.125 -6.22 12.295 -2.105 ;
      LAYER met1 ;
        RECT 3.39 -6.2 12.325 -5.91 ;
        RECT 11.94 -2.415 12.325 -2.125 ;
      LAYER mcon ;
        RECT 12.125 -2.355 12.295 -2.185 ;
        RECT 12.125 -6.14 12.295 -5.97 ;
    END
  END Vg_8
  PIN Vg_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.18 -6.77 13.35 -2.1 ;
      LAYER met1 ;
        RECT 3.445 -6.75 13.38 -6.46 ;
        RECT 12.94 -2.41 13.38 -2.12 ;
      LAYER mcon ;
        RECT 13.18 -2.35 13.35 -2.18 ;
        RECT 13.18 -6.69 13.35 -6.52 ;
    END
  END Vg_9
  PIN Vout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.6 1.285 23.08 14.235 ;
        RECT 22.67 1.285 22.93 14.27 ;
      LAYER li1 ;
        RECT 20.41 -1.87 20.58 1.185 ;
        RECT 20.395 10.48 20.565 13.405 ;
        RECT 19.355 -1.87 19.525 1.185 ;
        RECT 19.335 10.48 19.505 13.425 ;
        RECT 18.295 -1.87 18.465 1.185 ;
        RECT 18.275 10.48 18.445 13.42 ;
        RECT 16.62 -1.87 16.79 1.21 ;
        RECT 16.41 10.48 16.58 13.425 ;
        RECT 15.56 -1.87 15.73 1.21 ;
        RECT 15.35 10.48 15.52 13.425 ;
        RECT 14.5 -1.865 14.67 1.215 ;
        RECT 14.3 10.485 14.47 13.43 ;
        RECT 13.44 -1.865 13.61 1.215 ;
        RECT 13.245 10.485 13.415 13.43 ;
        RECT 12.385 -1.865 12.555 1.215 ;
        RECT 12.19 10.485 12.36 13.43 ;
        RECT 11.33 -1.865 11.5 1.215 ;
        RECT 11.13 10.485 11.3 13.42 ;
        RECT 9.715 -1.865 9.885 1.215 ;
        RECT 9.275 10.485 9.445 13.43 ;
        RECT 8.655 -1.865 8.825 1.215 ;
        RECT 8.22 10.485 8.39 13.43 ;
        RECT 7.595 -1.865 7.765 1.215 ;
        RECT 7.165 10.485 7.335 13.43 ;
        RECT 6.535 -1.865 6.705 1.215 ;
        RECT 6.105 10.485 6.275 13.43 ;
        RECT 5.48 -1.865 5.65 1.215 ;
        RECT 5.045 10.485 5.215 13.425 ;
        RECT 4.42 -1.865 4.59 1.22 ;
        RECT 3.985 10.485 4.155 13.44 ;
        RECT 3.36 -1.865 3.53 1.21 ;
        RECT 2.925 10.485 3.095 13.425 ;
      LAYER met1 ;
        RECT 2.165 1.45 23.06 2.07 ;
        RECT 22.735 1.425 22.995 2.07 ;
        RECT 20.38 0.875 20.61 2.07 ;
        RECT 19.325 0.875 19.555 2.07 ;
        RECT 18.265 0.875 18.495 2.07 ;
        RECT 16.59 0.9 16.82 2.07 ;
        RECT 15.53 0.9 15.76 2.07 ;
        RECT 14.47 0.905 14.7 2.07 ;
        RECT 13.41 0.905 13.64 2.07 ;
        RECT 12.355 0.905 12.585 2.07 ;
        RECT 11.3 0.905 11.53 2.07 ;
        RECT 9.685 0.905 9.915 2.07 ;
        RECT 8.625 0.905 8.855 2.07 ;
        RECT 7.565 0.905 7.795 2.07 ;
        RECT 6.505 0.905 6.735 2.07 ;
        RECT 5.45 0.905 5.68 2.07 ;
        RECT 4.39 0.91 4.62 2.07 ;
        RECT 3.33 0.9 3.56 2.07 ;
        RECT 2.045 13.64 23.035 14.29 ;
        RECT 22.67 13.63 22.93 14.29 ;
        RECT 20.365 13.095 20.595 14.29 ;
        RECT 19.305 13.115 19.535 14.29 ;
        RECT 18.245 13.11 18.475 14.29 ;
        RECT 16.38 13.115 16.61 14.29 ;
        RECT 15.32 13.115 15.55 14.29 ;
        RECT 14.27 13.12 14.5 14.29 ;
        RECT 13.215 13.12 13.445 14.29 ;
        RECT 12.16 13.12 12.39 14.29 ;
        RECT 11.1 13.11 11.33 14.29 ;
        RECT 9.245 13.12 9.475 14.29 ;
        RECT 8.19 13.12 8.42 14.29 ;
        RECT 7.135 13.12 7.365 14.29 ;
        RECT 6.075 13.12 6.305 14.29 ;
        RECT 5.015 13.115 5.245 14.29 ;
        RECT 3.955 13.13 4.185 14.29 ;
        RECT 2.895 13.115 3.125 14.29 ;
      LAYER mcon ;
        RECT 2.925 13.175 3.095 13.345 ;
        RECT 3.36 0.96 3.53 1.13 ;
        RECT 3.985 13.19 4.155 13.36 ;
        RECT 4.42 0.97 4.59 1.14 ;
        RECT 5.045 13.175 5.215 13.345 ;
        RECT 5.48 0.965 5.65 1.135 ;
        RECT 6.105 13.18 6.275 13.35 ;
        RECT 6.535 0.965 6.705 1.135 ;
        RECT 7.165 13.18 7.335 13.35 ;
        RECT 7.595 0.965 7.765 1.135 ;
        RECT 8.22 13.18 8.39 13.35 ;
        RECT 8.655 0.965 8.825 1.135 ;
        RECT 9.275 13.18 9.445 13.35 ;
        RECT 9.715 0.965 9.885 1.135 ;
        RECT 11.13 13.17 11.3 13.34 ;
        RECT 11.33 0.965 11.5 1.135 ;
        RECT 12.19 13.18 12.36 13.35 ;
        RECT 12.385 0.965 12.555 1.135 ;
        RECT 13.245 13.18 13.415 13.35 ;
        RECT 13.44 0.965 13.61 1.135 ;
        RECT 14.3 13.18 14.47 13.35 ;
        RECT 14.5 0.965 14.67 1.135 ;
        RECT 15.35 13.175 15.52 13.345 ;
        RECT 15.56 0.96 15.73 1.13 ;
        RECT 16.41 13.175 16.58 13.345 ;
        RECT 16.62 0.96 16.79 1.13 ;
        RECT 18.275 13.17 18.445 13.34 ;
        RECT 18.295 0.935 18.465 1.105 ;
        RECT 19.335 13.175 19.505 13.345 ;
        RECT 19.355 0.935 19.525 1.105 ;
        RECT 20.395 13.155 20.565 13.325 ;
        RECT 20.41 0.935 20.58 1.105 ;
      LAYER via ;
        RECT 22.725 14.035 22.875 14.185 ;
        RECT 22.725 13.715 22.875 13.865 ;
        RECT 22.79 1.83 22.94 1.98 ;
        RECT 22.79 1.51 22.94 1.66 ;
    END
  END Vout
END pass_transistors

END LIBRARY
