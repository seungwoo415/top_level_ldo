*.include "/home/ff/eecs251b/sky130/sky130_cds/sky130_release_0.0.1/models/sky130.lib.spice" section=tt
*.include "/home/ff/eecs251b/sky130/sky130_cds/sky130_release_0.0.1/models/sky130.lib.spice" tt


.SUBCKT pass_transistors Vg_0 Vg_1 Vg_2 Vg_3 Vg_4 Vg_5 Vg_6 Vg_7 Vg_8 Vg_9 Vg_10 Vg_11 Vg_12 Vg_13 Vg_14 Vg_15 Vg_16 Vg_17 Vg_18 Vg_19 Vg_20 Vg_21 Vg_22 Vg_23 Vg_24 Vg_25 Vg_26 Vg_27 Vg_28 Vg_29 Vg_30 Vg_31 Vout VDD 
 
   M1 Vout Vg_0 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M2 Vout Vg_1 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M3 Vout Vg_2 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M4 Vout Vg_3 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M5 Vout Vg_4 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M6 Vout Vg_5 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M7 Vout Vg_6 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M8 Vout Vg_7 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M9 Vout Vg_8 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M10 Vout Vg_9 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M11 Vout Vg_10 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M12 Vout Vg_11 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M13 Vout Vg_12 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M14 Vout Vg_13 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M15 Vout Vg_14 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M16 Vout Vg_15 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M17 Vout Vg_16 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M18 Vout Vg_17 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M19 Vout Vg_18 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M20 Vout Vg_19 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M21 Vout Vg_20 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M22 Vout Vg_21 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M23 Vout Vg_22 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M24 Vout Vg_23 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M25 Vout Vg_24 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M26 Vout Vg_25 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M27 Vout Vg_26 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M28 Vout Vg_27 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M29 Vout Vg_28 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M30 Vout Vg_29 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M31 Vout Vg_30 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
   M32 Vout Vg_31 VDD VDD pfet_01v8 l=0.25u nf=1 w=1.2u
.ENDS pass_transistors
