*
*
*
*                       LINUX           Wed Oct 30 02:49:35 2024
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 22.1.1-p041
*  Build Date     : Mon Apr 17 07:36:05 PDT 2023
*
*  HSPICE LIBRARY
*
*  OPERATING_TEMPERATURE 25
*  QRC_TECH_DIR /home/ff/eecs251b/sky130/sky130_cds/sky130_release_0.0.1/quantus/extraction/typical 
*
*
*

*
.SUBCKT pass_transistors Vg_22 Vg_12 Vg_29 Vg_16 Vg_6 Vg_23 Vg_13 Vg_0 Vg_17
+ Vg_7 Vg_30 Vg_24 Vg_14 Vg_1 Vg_8 Vg_18 Vg_31 Vg_25 Vg_15 Vg_2 Vg_9 Vg_19 VDD
+ Vg_3 Vg_26 Vout Vg_10 Vg_20 Vg_4 Vg_27 Vg_11 Vg_21 Vg_5 Vg_28
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MX159/X1/M0	Vout#118	Vg_14#1	VDD#130	VDD
+ pfet_01v8	L=2.5e-07	W=1.2e-06
MX159/X0/M0	Vout#110	Vg_13#1	VDD#122	VDD
+ pfet_01v8	L=2.5e-07	W=1.2e-06
MX158/X1/M0	Vout#114	Vg_30#1	VDD#126	VDD
+ pfet_01v8	L=2.5e-07	W=1.2e-06
MX158/X0/M0	Vout#106	Vg_29#1	VDD#118	VDD
+ pfet_01v8	L=2.5e-07	W=1.2e-06
MX157/X1/M0	Vout#102	Vg_12#1	VDD#110	VDD
+ pfet_01v8	L=2.5e-07	W=1.2e-06
MX157/X0/M0	Vout#94	Vg_11#1	VDD#102	VDD
+ pfet_01v8	L=2.5e-07	W=1.2e-06
MX156/X1/M0	Vout#98	Vg_28#1	VDD#106	VDD
+ pfet_01v8	L=2.5e-07	W=1.2e-06
MX156/X0/M0	Vout#90	Vg_27#1	VDD#98	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX155/X1/M0	Vout#86	Vg_10#1	VDD#94	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX155/X0/M0	Vout#78	Vg_9#1	VDD#86	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX154/X1/M0	Vout#66	Vg_24#1	VDD#74	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX154/X0/M0	Vout#58	Vg_23#1	VDD#66	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX153/X1/M0	Vout#46	Vg_5#1	VDD#50	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX153/X0/M0	Vout#38	Vg_4#1	VDD#42	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX152/X1/M0	Vout#26	Vg_19#1	VDD#30	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX152/X0/M0	Vout#18	Vg_18#1	VDD#22	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX151/X1/M0	Vout#14	Vg_1#1	VDD#18	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX151/X0/M0	Vout#6	Vg_0#1	VDD#10	VDD	pfet_01v8	L=2.5e-07
+ W=1.2e-06
MX150/X1/M0	Vout#10	Vg_17#1	VDD#14	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX150/X0/M0	Vout#2	Vg_16#1	VDD#6	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX149/M0	Vout#126	Vg_15#1	VDD#138	VDD
+ pfet_01v8	L=2.5e-07	W=1.2e-06
MX148/M0	Vout#122	Vg_31#1	VDD#134	VDD
+ pfet_01v8	L=2.5e-07	W=1.2e-06
MX147/M0	Vout#82	Vg_26#1	VDD#90	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX146/M0	Vout#74	Vg_25#1	VDD#82	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX145/M0	Vout#70	Vg_8#1	VDD#78	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX144/M0	Vout#62	Vg_7#1	VDD#70	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX143/M0	Vout#54	Vg_6#1	VDD#58	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX142/M0	Vout#50	Vg_22#1	VDD#54	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX141/M0	Vout#42	Vg_21#1	VDD#46	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX140/M0	Vout#34	Vg_20#1	VDD#38	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX139/M0	Vout#30	Vg_3#1	VDD#34	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
MX138/M0	Vout#22	Vg_2#1	VDD#26	VDD	pfet_01v8
+ L=2.5e-07	W=1.2e-06
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rg1	Vg_16#1	Vg_16#3	195.434387	$poly
Rg2	Vg_0#1	Vg_0#3	196.398376	$poly
Rg3	Vg_17#1	Vg_17#3	197.191559	$poly
Rg4	Vg_1#1	Vg_1#3	192.542389	$poly
Rg5	Vg_18#1	Vg_18#3	195.263565	$poly
Rg6	Vg_2#1	Vg_2#3	190.443558	$poly
Rg7	Vg_19#1	Vg_19#3	194.299561	$poly
Rg8	Vg_3#1	Vg_3#3	191.578384	$poly
Rg9	Vg_20#1	Vg_20#3	193.506378	$poly
Rg10	Vg_4#1	Vg_4#3	192.542389	$poly
Rg11	Vg_21#1	Vg_21#3	193.335556	$poly
Rg12	Vg_5#1	Vg_5#3	192.371567	$poly
Rg13	Vg_22#1	Vg_22#3	193.335556	$poly
Rg14	Vg_6#1	Vg_6#3	194.299561	$poly
Rg15	Vg_23#1	Vg_23#3	194.470383	$poly
Rg16	Vg_7#1	Vg_7#3	194.299561	$poly
Rg17	Vg_24#1	Vg_24#3	192.542389	$poly
Rg18	Vg_8#1	Vg_8#3	191.407562	$poly
Rg19	Vg_25#1	Vg_25#3	192.371567	$poly
Rg20	Vg_9#1	Vg_9#3	190.443558	$poly
Rg21	Vg_26#1	Vg_26#3	189.479553	$poly
Rg22	Vg_10#1	Vg_10#3	190.614380	$poly
Rg23	Vg_27#1	Vg_27#3	190.443558	$poly
Rg24	Vg_11#1	Vg_11#3	191.578384	$poly
Rg25	Vg_28#1	Vg_28#3	190.614380	$poly
Rg26	Vg_12#1	Vg_12#3	190.443558	$poly
Rg27	Vg_29#1	Vg_29#3	188.515564	$poly
Rg28	Vg_13#1	Vg_13#3	195.434387	$poly
Rg29	Vg_30#1	Vg_30#3	190.614380	$poly
Rg30	Vg_14#1	Vg_14#3	193.506378	$poly
Rg31	Vg_31#1	Vg_31#3	190.443558	$poly
Rg32	Vg_15#1	Vg_15#3	194.299561	$poly
Rf3	VDD#5	VDD#7	73.411766	$li
Rf5	VDD#6	VDD#7	5.000000	$li
Rf6	Vg_16#4	Vg_16#3	15.000000	$li
Rf7	VDD#9	VDD#11	76.047058	$li
Rf9	VDD#10	VDD#11	5.000000	$li
Rf10	Vout#1	Vout#3	163.764709	$li
Rf12	Vout#2	Vout#3	5.000000	$li
Rf13	Vg_0#4	Vg_0#3	15.000000	$li
Rf14	Vout#5	Vout#7	173.929413	$li
Rf16	Vout#6	Vout#7	5.000000	$li
Rf17	VDD#13	VDD#15	73.788239	$li
Rf19	VDD#14	VDD#15	5.000000	$li
Rf20	Vg_17#4	Vg_17#3	15.000000	$li
Rf22	VDD#17	VDD#19	76.047058	$li
Rf24	VDD#18	VDD#19	5.000000	$li
Rf25	Vout#9	Vout#11	164.894119	$li
Rf27	Vout#10	Vout#11	5.000000	$li
Rf28	Vg_1#4	Vg_1#3	15.000000	$li
Rf30	Vout#13	Vout#15	174.682343	$li
Rf32	Vout#14	Vout#15	5.000000	$li
Rf33	VDD#21	VDD#23	73.788239	$li
Rf35	VDD#22	VDD#23	5.000000	$li
Rf36	Vg_18#4	Vg_18#3	15.000000	$li
Rf38	VDD#25	VDD#27	76.047058	$li
Rf40	VDD#26	VDD#27	5.000000	$li
Rf41	Vout#17	Vout#19	163.764709	$li
Rf43	Vout#18	Vout#19	5.000000	$li
Rf44	Vg_2#4	Vg_2#3	15.000000	$li
Rf46	Vout#21	Vout#23	174.305878	$li
Rf48	Vout#22	Vout#23	5.000000	$li
Rf49	VDD#29	VDD#31	74.917648	$li
Rf51	VDD#30	VDD#31	5.000000	$li
Rf52	Vg_19#4	Vg_19#3	15.000000	$li
Rf54	VDD#33	VDD#35	76.047058	$li
Rf56	VDD#34	VDD#35	5.000000	$li
Rf57	Vout#25	Vout#27	164.141174	$li
Rf59	Vout#26	Vout#27	5.000000	$li
Rf60	Vg_3#4	Vg_3#3	15.000000	$li
Rf62	Vout#29	Vout#31	174.305878	$li
Rf64	Vout#30	Vout#31	5.000000	$li
Rf65	VDD#37	VDD#39	74.917648	$li
Rf67	VDD#38	VDD#39	5.000000	$li
Rf68	Vg_20#4	Vg_20#3	15.000000	$li
Rf70	VDD#41	VDD#43	76.047058	$li
Rf72	VDD#42	VDD#43	5.000000	$li
Rf73	Vout#33	Vout#35	164.141174	$li
Rf75	Vout#34	Vout#35	5.000000	$li
Rf76	Vg_4#4	Vg_4#3	15.000000	$li
Rf78	Vout#37	Vout#39	174.305878	$li
Rf80	Vout#38	Vout#39	5.000000	$li
Rf81	VDD#45	VDD#47	75.294113	$li
Rf83	VDD#46	VDD#47	5.000000	$li
Rf84	Vg_21#4	Vg_21#3	15.000000	$li
Rf86	VDD#49	VDD#51	76.047058	$li
Rf88	VDD#50	VDD#51	5.000000	$li
Rf89	Vout#41	Vout#43	164.141174	$li
Rf91	Vout#42	Vout#43	5.000000	$li
Rf92	Vg_5#4	Vg_5#3	15.000000	$li
Rf94	Vout#45	Vout#47	174.305878	$li
Rf96	Vout#46	Vout#47	5.000000	$li
Rf97	VDD#53	VDD#55	75.294113	$li
Rf99	VDD#54	VDD#55	5.000000	$li
Rf100	Vg_22#4	Vg_22#3	15.000000	$li
Rf102	VDD#57	VDD#59	76.423531	$li
Rf104	VDD#58	VDD#59	5.000000	$li
Rf105	Vout#49	Vout#51	164.141174	$li
Rf107	Vout#50	Vout#51	5.000000	$li
Rf108	Vg_6#4	Vg_6#3	15.000000	$li
Rf110	Vout#53	Vout#55	174.305878	$li
Rf112	Vout#54	Vout#55	5.000000	$li
Rf115	VDD#65	VDD#67	74.541176	$li
Rf117	VDD#66	VDD#67	5.000000	$li
Rf118	VDD#69	VDD#71	76.047058	$li
Rf120	VDD#70	VDD#71	5.000000	$li
Rf121	Vg_23#4	Vg_23#3	15.000000	$li
Rf123	Vg_7#4	Vg_7#3	15.000000	$li
Rf125	Vout#57	Vout#59	163.388229	$li
Rf127	Vout#58	Vout#59	5.000000	$li
Rf128	Vout#61	Vout#63	174.305878	$li
Rf130	Vout#62	Vout#63	5.000000	$li
Rf131	VDD#73	VDD#75	74.541176	$li
Rf133	VDD#74	VDD#75	5.000000	$li
Rf134	VDD#77	VDD#79	76.047058	$li
Rf136	VDD#78	VDD#79	5.000000	$li
Rf137	Vg_24#4	Vg_24#3	15.000000	$li
Rf139	Vg_8#4	Vg_8#3	15.000000	$li
Rf141	Vout#65	Vout#67	164.141174	$li
Rf143	Vout#66	Vout#67	5.000000	$li
Rf144	Vout#69	Vout#71	174.305878	$li
Rf146	Vout#70	Vout#71	5.000000	$li
Rf147	VDD#81	VDD#83	74.541176	$li
Rf149	VDD#82	VDD#83	5.000000	$li
Rf150	VDD#85	VDD#87	76.047058	$li
Rf152	VDD#86	VDD#87	5.000000	$li
Rf153	Vg_25#4	Vg_25#3	15.000000	$li
Rf155	Vg_9#4	Vg_9#3	15.000000	$li
Rf157	Vout#73	Vout#75	164.141174	$li
Rf159	Vout#74	Vout#75	5.000000	$li
Rf160	Vout#77	Vout#79	174.305878	$li
Rf162	Vout#78	Vout#79	5.000000	$li
Rf163	VDD#89	VDD#91	74.541176	$li
Rf165	VDD#90	VDD#91	5.000000	$li
Rf166	VDD#93	VDD#95	76.047058	$li
Rf168	VDD#94	VDD#95	5.000000	$li
Rf169	Vg_26#4	Vg_26#3	15.000000	$li
Rf171	Vg_10#4	Vg_10#3	15.000000	$li
Rf173	Vout#81	Vout#83	164.141174	$li
Rf175	Vout#82	Vout#83	5.000000	$li
Rf176	Vout#85	Vout#87	174.305878	$li
Rf178	Vout#86	Vout#87	5.000000	$li
Rf179	VDD#97	VDD#99	74.164703	$li
Rf181	VDD#98	VDD#99	5.000000	$li
Rf182	VDD#101	VDD#103	76.047058	$li
Rf184	VDD#102	VDD#103	5.000000	$li
Rf185	Vg_27#4	Vg_27#3	15.000000	$li
Rf187	Vg_11#4	Vg_11#3	15.000000	$li
Rf189	Vout#89	Vout#91	164.141174	$li
Rf191	Vout#90	Vout#91	5.000000	$li
Rf192	Vout#93	Vout#95	174.305878	$li
Rf194	Vout#94	Vout#95	5.000000	$li
Rf195	VDD#105	VDD#107	74.917648	$li
Rf197	VDD#106	VDD#107	5.000000	$li
Rf198	VDD#109	VDD#111	76.047058	$li
Rf200	VDD#110	VDD#111	5.000000	$li
Rf201	Vg_28#4	Vg_28#3	15.000000	$li
Rf203	Vg_12#4	Vg_12#3	15.000000	$li
Rf205	Vout#97	Vout#99	164.141174	$li
Rf207	Vout#98	Vout#99	5.000000	$li
Rf208	Vout#101	Vout#103	174.305878	$li
Rf210	Vout#102	Vout#103	5.000000	$li
Rf213	VDD#117	VDD#119	74.917648	$li
Rf215	VDD#118	VDD#119	5.000000	$li
Rf216	VDD#121	VDD#123	76.047058	$li
Rf218	VDD#122	VDD#123	5.000000	$li
Rf219	Vg_29#4	Vg_29#3	15.000000	$li
Rf221	Vg_13#4	Vg_13#3	15.000000	$li
Rf223	Vout#105	Vout#107	163.764709	$li
Rf225	Vout#106	Vout#107	5.000000	$li
Rf226	Vout#109	Vout#111	172.423538	$li
Rf228	Vout#110	Vout#111	5.000000	$li
Rf229	VDD#125	VDD#127	76.423531	$li
Rf231	VDD#126	VDD#127	5.000000	$li
Rf232	VDD#129	VDD#131	76.047058	$li
Rf234	VDD#130	VDD#131	5.000000	$li
Rf235	Vg_30#4	Vg_30#3	15.000000	$li
Rf237	Vg_14#4	Vg_14#3	15.000000	$li
Rf239	Vout#113	Vout#115	164.141174	$li
Rf241	Vout#114	Vout#115	5.000000	$li
Rf242	Vout#117	Vout#119	172.423538	$li
Rf244	Vout#118	Vout#119	5.000000	$li
Rf245	VDD#133	VDD#135	75.294113	$li
Rf247	VDD#134	VDD#135	5.000000	$li
Rf248	VDD#137	VDD#139	76.047058	$li
Rf250	VDD#138	VDD#139	5.000000	$li
Rf251	Vg_31#4	Vg_31#3	15.000000	$li
Rf253	Vg_15#4	Vg_15#3	15.000000	$li
Rf255	Vout#121	Vout#123	162.635284	$li
Rf257	Vout#122	Vout#123	5.000000	$li
Rf258	Vout#125	Vout#127	172.423538	$li
Rf260	Vout#126	Vout#127	5.000000	$li
Re1	Vg_16#4	Vg_16	152.002151	$metal1
Re2	Vg_0#6	Vg_0#4	152.005737	$metal1
Re3	Vg_0	Vg_0#8	0.005740	$metal1
Re4	Vg_0#6	Vg_0#8	0.034483	$metal1
Re5	Vg_17#4	Vg_17	152.009033	$metal1
Re6	Vg_1#7	Vg_1#4	152.006531	$metal1
Re7	Vg_1	Vg_1#9	0.006530	$metal1
Re8	Vg_1#7	Vg_1#9	0.021552	$metal1
Re9	Vg_18	Vg_18#4	152.010773	$metal1
Re10	Vg_2#4	Vg_2	152.004303	$metal1
Re11	Vg_19#4	Vg_19	152.002151	$metal1
Re12	Vg_3	Vg_3#4	152.007721	$metal1
Re13	Vg_20#4	Vg_20	152.004303	$metal1
Re14	Vg_4	Vg_4#4	152.002151	$metal1
Re15	Vg_21	Vg_21#4	152.006470	$metal1
Re16	Vg_5	Vg_5#4	152.002151	$metal1
Re17	Vg_22	Vg_22#4	152.005142	$metal1
Re18	Vg_6	Vg_6#4	152.004303	$metal1
Re19	Vg_23#4	Vg_23	152.006470	$metal1
Re20	Vg_7	Vg_7#4	152.008453	$metal1
Re21	Vg_24	Vg_24#4	152.009506	$metal1
Re22	Vg_8#4	Vg_8	152.010773	$metal1
Re23	Vg_25	Vg_25#4	152.010773	$metal1
Re24	Vg_9#4	Vg_9	152.004257	$metal1
Re25	Vg_26	Vg_26#4	152.015091	$metal1
Re26	Vg_10#4	Vg_10	152.004074	$metal1
Re27	Vg_27	Vg_27#4	152.006470	$metal1
Re28	Vg_11	Vg_11#4	152.008621	$metal1
Re29	Vg_28	Vg_28#4	152.021545	$metal1
Re30	Vg_12	Vg_12#4	152.007629	$metal1
Re31	Vg_29#4	Vg_29	152.012924	$metal1
Re32	Vg_13	Vg_13#4	152.002151	$metal1
Re33	Vg_30#7	Vg_30	0.005000	$metal1
Re34	Vg_30#4	Vg_30#9	152.005005	$metal1
Re35	Vg_30#7	Vg_30#9	0.023707	$metal1
Re36	Vg_14#4	Vg_14	152.017242	$metal1
Re37	Vg_31	Vg_31#4	152.012924	$metal1
Re38	Vg_15	Vg_15#4	152.002808	$metal1
Re41	VDD#147	VDD#148	0.241701	$metal1
Re42	VDD#148	VDD#149	0.242858	$metal1
Re43	VDD#149	VDD#150	0.124803	$metal1
Re44	VDD#150	VDD#151	0.257904	$metal1
Re45	VDD#151	VDD#152	0.242858	$metal1
Re46	VDD#152	VDD#153	0.242858	$metal1
Re47	VDD#153	VDD#154	0.242858	$metal1
Re48	VDD#154	VDD#155	0.241701	$metal1
Re49	VDD#155	VDD#156	0.241701	$metal1
Re50	VDD#156	VDD#157	0.112071	$metal1
Re51	VDD#157	VDD#158	0.256747	$metal1
Re52	VDD#158	VDD#159	0.242858	$metal1
Re53	VDD#159	VDD#160	0.242858	$metal1
Re54	VDD#160	VDD#161	0.242858	$metal1
Re55	VDD#161	VDD#162	0.241701	$metal1
Re56	VDD#162	VDD#163	0.242858	$metal1
Re57	VDD#163	VDD#164	0.242858	$metal1
Re58	VDD#164	VDD#3	0.170040	$metal1
Re59	VDD#3	VDD#166	0.385344	$metal1
Re60	VDD#147	VDD#137	152.211960	$metal1
Re61	VDD#148	VDD#129	152.211960	$metal1
Re62	VDD#149	VDD#121	152.211960	$metal1
Re64	VDD#151	VDD#109	152.211960	$metal1
Re65	VDD#152	VDD#101	152.211960	$metal1
Re66	VDD#153	VDD#93	152.209244	$metal1
Re67	VDD#154	VDD#85	152.209244	$metal1
Re68	VDD#155	VDD#77	152.209244	$metal1
Re69	VDD#156	VDD#69	152.209244	$metal1
Re71	VDD#158	VDD#57	152.206528	$metal1
Re72	VDD#159	VDD#49	152.209244	$metal1
Re73	VDD#160	VDD#41	152.209244	$metal1
Re74	VDD#161	VDD#33	152.209244	$metal1
Re75	VDD#162	VDD#25	152.209244	$metal1
Re76	VDD#163	VDD#17	152.209244	$metal1
Re77	VDD#164	VDD#9	152.209244	$metal1
Re78	VDD	VDD#141	0.224537	$metal1
Re79	VDD#141	VDD#186	0.277679	$metal1
Re80	VDD#186	VDD#187	0.242858	$metal1
Re81	VDD#187	VDD#188	0.242858	$metal1
Re82	VDD#188	VDD#189	0.150266	$metal1
Re83	VDD#189	VDD#190	0.276423	$metal1
Re84	VDD#190	VDD#191	0.242858	$metal1
Re85	VDD#191	VDD#192	0.240543	$metal1
Re86	VDD#192	VDD#193	0.241701	$metal1
Re87	VDD#193	VDD#194	0.241701	$metal1
Re88	VDD#194	VDD#195	0.242858	$metal1
Re89	VDD#195	VDD#196	0.151423	$metal1
Re90	VDD#196	VDD#197	0.272951	$metal1
Re91	VDD#197	VDD#198	0.241701	$metal1
Re92	VDD#198	VDD#199	0.241701	$metal1
Re93	VDD#199	VDD#200	0.242858	$metal1
Re94	VDD#200	VDD#201	0.242858	$metal1
Re95	VDD#201	VDD#202	0.242858	$metal1
Re96	VDD#202	VDD#203	0.242858	$metal1
Re97	VDD#203	VDD#1	0.160781	$metal1
Re98	VDD#1	VDD#205	0.296467	$metal1
Re99	VDD#186	VDD#133	152.217392	$metal1
Re100	VDD#187	VDD#125	152.209244	$metal1
Re101	VDD#188	VDD#117	152.220108	$metal1
Re103	VDD#190	VDD#105	152.220108	$metal1
Re104	VDD#191	VDD#97	152.225540	$metal1
Re105	VDD#192	VDD#89	152.220108	$metal1
Re106	VDD#193	VDD#81	152.220108	$metal1
Re107	VDD#194	VDD#73	152.220108	$metal1
Re108	VDD#195	VDD#65	152.220108	$metal1
Re110	VDD#197	VDD#53	152.214676	$metal1
Re111	VDD#198	VDD#45	152.214676	$metal1
Re112	VDD#199	VDD#37	152.217392	$metal1
Re113	VDD#200	VDD#29	152.217392	$metal1
Re114	VDD#201	VDD#21	152.225540	$metal1
Re115	VDD#202	VDD#13	152.225540	$metal1
Re116	VDD#203	VDD#5	152.228256	$metal1
Re117	Vout#121	Vout#130	152.270981	$metal1
Re118	Vout#130	Vout#131	0.202016	$metal1
Re119	Vout#131	Vout#132	0.202016	$metal1
Re120	Vout#132	Vout#133	0.356823	$metal1
Re121	Vout#133	Vout#134	0.202016	$metal1
Re122	Vout#134	Vout#135	0.200093	$metal1
Re123	Vout#135	Vout#136	0.201054	$metal1
Re124	Vout#136	Vout#137	0.201054	$metal1
Re125	Vout#137	Vout#138	0.202016	$metal1
Re126	Vout#138	Vout#139	0.354900	$metal1
Re127	Vout#139	Vout#140	0.201054	$metal1
Re128	Vout#140	Vout#141	0.201054	$metal1
Re129	Vout#141	Vout#142	0.202016	$metal1
Re130	Vout#142	Vout#143	0.202016	$metal1
Re131	Vout#143	Vout#144	0.202016	$metal1
Re132	Vout#144	Vout#1	152.462936	$metal1
Re133	Vout#130	Vout	0.299085	$metal1
Re134	Vout	Vout#146	0.145803	$metal1
Re135	Vout#131	Vout#113	152.260117	$metal1
Re136	Vout#132	Vout#105	152.262833	$metal1
Re137	Vout#133	Vout#97	152.260117	$metal1
Re138	Vout#134	Vout#89	152.260117	$metal1
Re139	Vout#135	Vout#81	152.257401	$metal1
Re140	Vout#136	Vout#73	152.257401	$metal1
Re141	Vout#137	Vout#65	152.257401	$metal1
Re142	Vout#138	Vout#57	152.262833	$metal1
Re143	Vout#139	Vout#49	152.257401	$metal1
Re144	Vout#140	Vout#41	152.257401	$metal1
Re145	Vout#141	Vout#33	152.257401	$metal1
Re146	Vout#142	Vout#25	152.257401	$metal1
Re147	Vout#143	Vout#17	152.260117	$metal1
Re148	Vout#144	Vout#9	152.251953	$metal1
Re149	Vout#125	Vout#162	152.285400	$metal1
Re150	Vout#162	Vout#163	0.210716	$metal1
Re151	Vout#163	Vout#164	0.211724	$metal1
Re152	Vout#164	Vout#165	0.335716	$metal1
Re153	Vout#165	Vout#166	0.211724	$metal1
Re154	Vout#166	Vout#167	0.211724	$metal1
Re155	Vout#167	Vout#168	0.211724	$metal1
Re156	Vout#168	Vout#169	0.210716	$metal1
Re157	Vout#169	Vout#170	0.210716	$metal1
Re158	Vout#170	Vout#171	0.323619	$metal1
Re159	Vout#171	Vout#172	0.211724	$metal1
Re160	Vout#172	Vout#173	0.211724	$metal1
Re161	Vout#173	Vout#174	0.211724	$metal1
Re162	Vout#174	Vout#175	0.210716	$metal1
Re163	Vout#175	Vout#176	0.211724	$metal1
Re164	Vout#176	Vout#177	0.211724	$metal1
Re166	Vout#162	Vout#179	0.475952	$metal1
Re167	Vout#163	Vout#117	152.285400	$metal1
Re168	Vout#164	Vout#109	152.285400	$metal1
Re169	Vout#165	Vout#101	152.271820	$metal1
Re170	Vout#166	Vout#93	152.271820	$metal1
Re171	Vout#167	Vout#85	152.269104	$metal1
Re172	Vout#168	Vout#77	152.269104	$metal1
Re173	Vout#169	Vout#69	152.269104	$metal1
Re174	Vout#170	Vout#61	152.269104	$metal1
Re175	Vout#171	Vout#53	152.269104	$metal1
Re176	Vout#172	Vout#45	152.269104	$metal1
Re177	Vout#173	Vout#37	152.269104	$metal1
Re178	Vout#174	Vout#29	152.269104	$metal1
Re179	Vout#175	Vout#21	152.269104	$metal1
Re180	Vout#176	Vout#13	152.266388	$metal1
Re181	Vout#177	Vout#5	152.271820	$metal1
Rd1	VDD#166	VDD#205	8.779514	$metal2
Rd2	Vout#179	Vout#146	7.678386	$metal2
*
*       CAPACITOR CARDS
*
*
C1	Vg_22	35	1.67999e-15
C2	Vg_12	35	2.64876e-15
C3	Vg_29	35	3.32448e-15
C4	Vg_16	35	1.3278e-16
C5	Vg_6	35	1.64602e-15
C6	Vg_23	35	1.83919e-15
C7	Vg_13	35	3.16762e-15
C8	Vg_17	35	4.05973e-16
C9	Vg_7	35	1.85173e-15
C10	Vg_30	35	3.85144e-15
C11	Vg_24	35	1.98457e-15
C12	Vg_14	35	3.9048e-15
C13	Vg_1	35	3.91524e-16
C14	Vg_8	35	2.00249e-15
C15	Vg_18	35	6.93037e-16
C16	Vg_31	35	3.36252e-15
C17	Vg_25	35	2.54342e-15
C18	Vg_15	35	2.96471e-15
C19	Vg_2	35	6.6071e-16
C20	Vg_9	35	2.48229e-15
C21	Vg_19	35	9.8597e-16
C22	VDD	35	1.10909e-15
C23	Vg_3	35	9.61771e-16
C24	Vg_26	35	2.78092e-15
C25	Vout	35	1.26656e-16
C26	Vg_10	35	2.71927e-15
C27	Vg_20	35	1.23666e-15
C28	Vg_4	35	1.25126e-15
C29	Vg_27	35	2.51976e-15
C30	Vg_11	35	2.55814e-15
C31	Vg_21	35	1.48665e-15
C32	Vg_5	35	1.46459e-15
C33	Vg_28	35	2.76453e-15
C34	Vg_15#1	35	9.38371e-17
C35	Vg_31#1	35	9.39616e-17
C36	Vg_14#1	35	8.97204e-17
C37	Vg_30#1	35	9.07559e-17
C38	Vg_13#1	35	9.35208e-17
C39	Vg_29#1	35	9.45117e-17
C40	Vg_12#1	35	9.43835e-17
C41	Vg_28#1	35	9.42209e-17
C42	Vg_11#1	35	8.99623e-17
C43	Vg_27#1	35	9.03416e-17
C44	Vg_10#1	35	9.05381e-17
C45	Vg_26#1	35	9.0937e-17
C46	Vg_9#1	35	8.96047e-17
C47	Vg_25#1	35	8.9794e-17
C48	Vg_8#1	35	8.96347e-17
C49	Vg_24#1	35	8.9757e-17
C50	Vg_7#1	35	9.15124e-17
C51	Vg_23#1	35	9.41921e-17
C52	Vg_6#1	35	8.52175e-17
C53	Vg_22#1	35	9.30757e-17
C54	Vg_5#1	35	8.57571e-17
C55	Vg_21#1	35	8.59637e-17
C56	Vg_4#1	35	8.91961e-17
C57	Vg_20#1	35	8.53255e-17
C58	Vg_3#1	35	9.24427e-17
C59	Vg_19#1	35	8.83795e-17
C60	Vg_2#1	35	9.33234e-17
C61	Vg_18#1	35	9.34393e-17
C62	Vg_1#1	35	9.60742e-17
C63	Vg_17#1	35	9.48116e-17
C64	Vg_0#1	35	1.02003e-16
C65	Vg_16#1	35	1.00426e-16
C66	Vout#179	35	6.74554e-16
C67	Vout#146	35	5.72488e-16
C68	VDD#166	35	6.36814e-16
C69	VDD#205	35	5.69281e-16
C70	VDD#141	35	1.65279e-16
C71	Vout#125	35	1.58608e-16
C72	Vout#121	35	1.77771e-16
C73	Vg_15#4	35	6.48836e-16
C74	Vg_31#4	35	6.53308e-16
C75	VDD#137	35	8.72651e-17
C76	VDD#133	35	9.48972e-17
C77	Vout#117	35	1.32682e-16
C78	Vout#113	35	1.46567e-16
C79	Vg_14#4	35	6.59781e-16
C80	Vg_30#4	35	6.61897e-16
C81	VDD#129	35	7.73647e-17
C82	VDD#125	35	7.92448e-17
C83	Vout#109	35	1.6256e-16
C84	Vout#105	35	1.75216e-16
C85	Vg_13#4	35	2.95691e-16
C86	Vg_29#4	35	2.96042e-16
C87	VDD#121	35	5.87429e-17
C88	VDD#117	35	6.15668e-17
C89	Vout#101	35	1.58836e-16
C90	Vout#97	35	1.7254e-16
C91	Vg_12#4	35	5.32275e-16
C92	Vg_28#4	35	5.27442e-16
C93	VDD#109	35	7.93141e-17
C94	VDD#105	35	8.23483e-17
C95	Vout#93	35	1.3336e-16
C96	Vout#89	35	1.47566e-16
C97	Vg_11#4	35	5.04787e-16
C98	Vg_27#4	35	5.03356e-16
C99	VDD#101	35	8.01937e-17
C100	VDD#97	35	8.03917e-17
C101	Vout#85	35	1.31089e-16
C102	Vout#81	35	1.44549e-16
C103	Vg_10#4	35	4.54706e-16
C104	Vg_26#4	35	4.60529e-16
C105	VDD#93	35	7.70329e-17
C106	VDD#89	35	7.95382e-17
C107	Vout#77	35	1.29354e-16
C108	Vout#73	35	1.43039e-16
C109	Vg_9#4	35	4.13623e-16
C110	Vg_25#4	35	4.12292e-16
C111	VDD#85	35	7.86639e-17
C112	VDD#81	35	8.08399e-17
C113	Vout#69	35	1.29417e-16
C114	Vout#65	35	1.44174e-16
C115	Vg_8#4	35	3.66684e-16
C116	Vg_24#4	35	3.63889e-16
C117	VDD#77	35	7.75144e-17
C118	VDD#73	35	8.03269e-17
C119	Vout#61	35	1.41983e-16
C120	Vout#57	35	1.75674e-16
C121	Vg_7#4	35	3.13066e-16
C122	Vg_23#4	35	3.11076e-16
C123	VDD#69	35	5.8526e-17
C124	VDD#65	35	6.06505e-17
C125	Vout#53	35	1.42056e-16
C126	Vg_6#4	35	2.66612e-16
C127	Vout#49	35	1.71665e-16
C128	VDD#57	35	7.72711e-17
C129	Vg_22#4	35	2.63702e-16
C130	VDD#53	35	8.33286e-17
C131	Vout#45	35	1.29576e-16
C132	Vg_5#4	35	2.3256e-16
C133	Vout#41	35	1.43735e-16
C134	VDD#49	35	8.00448e-17
C135	Vg_21#4	35	2.27345e-16
C136	VDD#45	35	7.99452e-17
C137	Vout#37	35	1.29687e-16
C138	Vg_4#4	35	1.88106e-16
C139	Vout#33	35	1.43387e-16
C140	VDD#41	35	7.82613e-17
C141	Vg_20#4	35	1.90181e-16
C142	VDD#37	35	8.22395e-17
C143	Vout#29	35	1.29497e-16
C144	Vg_3#4	35	1.53275e-16
C145	Vout#25	35	1.44758e-16
C146	VDD#33	35	7.85977e-17
C147	Vg_19#4	35	1.53972e-16
C148	VDD#29	35	7.93163e-17
C149	Vout#21	35	1.32172e-16
C150	Vg_2#4	35	1.14805e-16
C151	Vout#17	35	1.50154e-16
C152	VDD#25	35	7.83221e-17
C153	Vg_18#4	35	1.13959e-16
C154	VDD#21	35	7.78135e-17
C155	Vout#13	35	1.32311e-16
C156	Vg_1#4	35	7.30495e-17
C157	Vout#9	35	1.45023e-16
C158	VDD#17	35	7.82279e-17
C159	Vg_17#4	35	6.90543e-17
C160	VDD#13	35	7.4614e-17
C161	Vout#5	35	1.58616e-16
C162	Vg_0#4	35	4.34391e-17
C163	Vout#1	35	3.73517e-16
C164	VDD#9	35	6.88261e-17
C165	Vg_16#4	35	4.67908e-17
C166	VDD#5	35	6.67359e-17
C167	VDD#3	35	1.04876e-16
C168	VDD#1	35	4.51494e-17
C169	Vg_13#3	35	2.86649e-16
C170	Vg_29#3	35	2.85012e-16
C171	Vout#126	35	2.22217e-16
C172	Vout#122	35	1.90226e-16
C173	VDD#138	35	1.5516e-16
C174	VDD#134	35	1.54614e-16
C175	Vout#118	35	2.37542e-16
C176	Vout#114	35	2.24611e-16
C177	VDD#130	35	1.52548e-16
C178	VDD#126	35	1.53155e-16
C179	Vout#110	35	2.297e-16
C180	Vout#106	35	2.24325e-16
C181	VDD#122	35	9.59557e-17
C182	VDD#118	35	9.51442e-17
C183	Vout#102	35	2.26904e-16
C184	Vout#98	35	1.97911e-16
C185	VDD#110	35	1.48918e-16
C186	VDD#106	35	1.47503e-16
C187	Vout#94	35	2.49973e-16
C188	Vout#90	35	2.28655e-16
C189	VDD#102	35	1.56464e-16
C190	VDD#98	35	1.50945e-16
C191	Vout#86	35	2.4464e-16
C192	Vout#82	35	2.24379e-16
C193	VDD#94	35	1.55899e-16
C194	VDD#90	35	1.54752e-16
C195	Vout#78	35	2.44359e-16
C196	Vout#74	35	2.23132e-16
C197	VDD#86	35	1.55014e-16
C198	VDD#82	35	1.52507e-16
C199	Vout#70	35	2.45287e-16
C200	Vout#66	35	2.23426e-16
C201	VDD#78	35	1.47892e-16
C202	VDD#74	35	1.56233e-16
C203	Vout#62	35	2.39607e-16
C204	Vout#58	35	2.23915e-16
C205	VDD#70	35	9.51129e-17
C206	VDD#66	35	9.59272e-17
C207	Vout#54	35	2.27228e-16
C208	Vout#50	35	1.99129e-16
C209	VDD#58	35	1.46609e-16
C210	VDD#54	35	1.46142e-16
C211	Vout#46	35	2.48462e-16
C212	Vout#42	35	2.29936e-16
C213	VDD#50	35	1.50078e-16
C214	VDD#46	35	1.48095e-16
C215	Vout#38	35	2.43872e-16
C216	Vout#34	35	2.22588e-16
C217	VDD#42	35	1.52145e-16
C218	VDD#38	35	1.48631e-16
C219	Vout#30	35	2.44046e-16
C220	Vout#26	35	2.21875e-16
C221	VDD#34	35	1.55117e-16
C222	VDD#30	35	1.54183e-16
C223	Vout#22	35	2.4604e-16
C224	Vout#18	35	2.22618e-16
C225	VDD#26	35	1.57644e-16
C226	VDD#22	35	1.57132e-16
C227	Vout#14	35	2.42815e-16
C228	Vout#10	35	2.20032e-16
C229	VDD#18	35	1.58809e-16
C230	VDD#14	35	1.58937e-16
C231	Vout#6	35	2.49377e-16
C232	Vout#2	35	2.27134e-16
C233	VDD#10	35	1.05882e-16
C234	VDD#6	35	1.04564e-16
C235	Vg_0#6	35	1.0896e-16
C236	Vg_0#8	35	3.73528e-17
C237	Vg_1#7	35	2.74351e-17
C238	Vg_1#9	35	1.89281e-17
C239	Vg_30#9	35	2.13062e-17
C240	VDD#147	35	4.2628e-16
C241	VDD#148	35	1.68538e-16
C242	VDD#149	35	1.06886e-16
C243	VDD#150	35	1.89505e-16
C244	VDD#151	35	1.81632e-16
C245	VDD#152	35	1.74333e-16
C246	VDD#153	35	1.74116e-16
C247	VDD#154	35	1.74137e-16
C248	VDD#155	35	1.73562e-16
C249	VDD#157	35	2.8592e-16
C250	VDD#158	35	1.77973e-16
C251	VDD#159	35	1.74168e-16
C252	VDD#160	35	1.74938e-16
C253	VDD#161	35	1.73994e-16
C254	VDD#162	35	1.735e-16
C255	VDD#163	35	1.74326e-16
C256	VDD#164	35	1.14079e-16
C257	VDD#186	35	1.7707e-16
C258	VDD#187	35	1.80427e-16
C259	VDD#188	35	1.20498e-16
C260	VDD#189	35	1.88436e-16
C261	VDD#190	35	1.95453e-16
C262	VDD#191	35	1.80204e-16
C263	VDD#192	35	1.78587e-16
C264	VDD#193	35	1.79157e-16
C265	VDD#194	35	1.79986e-16
C266	VDD#195	35	1.20764e-16
C267	VDD#196	35	1.91494e-16
C268	VDD#197	35	1.92436e-16
C269	VDD#198	35	1.78769e-16
C270	VDD#199	35	1.78899e-16
C271	VDD#200	35	1.79955e-16
C272	VDD#201	35	1.79693e-16
C273	VDD#202	35	1.80165e-16
C274	VDD#203	35	1.19309e-16
C275	Vout#130	35	1.51763e-16
C276	Vout#131	35	1.11068e-16
C277	Vout#132	35	1.61842e-16
C278	Vout#133	35	1.60971e-16
C279	Vout#134	35	1.0991e-16
C280	Vout#135	35	1.09403e-16
C281	Vout#136	35	1.10125e-16
C282	Vout#137	35	1.10551e-16
C283	Vout#138	35	1.61319e-16
C284	Vout#139	35	1.59904e-16
C285	Vout#140	35	1.10241e-16
C286	Vout#141	35	1.10432e-16
C287	Vout#142	35	1.1074e-16
C288	Vout#143	35	1.1038e-16
C289	Vout#144	35	1.25721e-16
C290	Vout#162	35	2.06854e-16
C291	Vout#163	35	1.41406e-16
C292	Vout#164	35	1.87215e-16
C293	Vout#165	35	1.85708e-16
C294	Vout#166	35	1.39798e-16
C295	Vout#167	35	1.39602e-16
C296	Vout#168	35	1.39231e-16
C297	Vout#169	35	1.38868e-16
C298	Vout#170	35	1.80358e-16
C299	Vout#171	35	1.79274e-16
C300	Vout#172	35	1.39607e-16
C301	Vout#173	35	1.39605e-16
C302	Vout#174	35	1.39231e-16
C303	Vout#175	35	1.39206e-16
C304	Vout#176	35	1.39645e-16
C305	Vout#177	35	2.59484e-16
*
*
.ENDS pass_transistors
*
